module controller_test; 

  localparam integer HLT=0, SKZ=1, ADD=2, AND=3, XOR=4, LDA=5, STO=6, JMP=7;

  reg [
  reg [

  wire [4:0] check_guess ; //wire for the check guess states 
  wire        win; //wire for winning  
  wire        lose; //wire for losing 

  
  controller controller_inst \


    
    
  
