VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 69.440 200.000 70.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 442.400 200.000 442.960 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 815.360 200.000 815.920 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 1188.320 200.000 1188.880 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 1561.280 200.000 1561.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 1934.240 200.000 1934.800 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 2307.200 200.000 2307.760 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 2680.160 200.000 2680.720 ;
    END
  END io_in[7]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 318.080 200.000 318.640 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1966.720 4.000 1967.280 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1592.640 4.000 1593.200 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1218.560 4.000 1219.120 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 844.480 4.000 845.040 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 470.400 4.000 470.960 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.320 4.000 96.880 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 691.040 200.000 691.600 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 1064.000 200.000 1064.560 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 1436.960 200.000 1437.520 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 1809.920 200.000 1810.480 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 2182.880 200.000 2183.440 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 2555.840 200.000 2556.400 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 2928.800 200.000 2929.360 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2714.880 4.000 2715.440 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2340.800 4.000 2341.360 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 193.760 200.000 194.320 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2153.760 4.000 2154.320 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1779.680 4.000 1780.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1405.600 4.000 1406.160 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1031.520 4.000 1032.080 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 657.440 4.000 658.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 283.360 4.000 283.920 ;
    END
  END io_out[15]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 566.720 200.000 567.280 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 939.680 200.000 940.240 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 1312.640 200.000 1313.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 1685.600 200.000 1686.160 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 2058.560 200.000 2059.120 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 2431.520 200.000 2432.080 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 2804.480 200.000 2805.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2901.920 4.000 2902.480 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2527.840 4.000 2528.400 ;
    END
  END io_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 2983.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 2983.420 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 2983.420 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 193.200 2983.420 ;
      LAYER Metal2 ;
        RECT 8.540 4.300 194.180 2983.310 ;
        RECT 8.540 4.000 48.980 4.300 ;
        RECT 50.140 4.000 148.660 4.300 ;
        RECT 149.820 4.000 194.180 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 2929.660 196.000 2983.260 ;
        RECT 4.000 2928.500 195.700 2929.660 ;
        RECT 4.000 2902.780 196.000 2928.500 ;
        RECT 4.300 2901.620 196.000 2902.780 ;
        RECT 4.000 2805.340 196.000 2901.620 ;
        RECT 4.000 2804.180 195.700 2805.340 ;
        RECT 4.000 2715.740 196.000 2804.180 ;
        RECT 4.300 2714.580 196.000 2715.740 ;
        RECT 4.000 2681.020 196.000 2714.580 ;
        RECT 4.000 2679.860 195.700 2681.020 ;
        RECT 4.000 2556.700 196.000 2679.860 ;
        RECT 4.000 2555.540 195.700 2556.700 ;
        RECT 4.000 2528.700 196.000 2555.540 ;
        RECT 4.300 2527.540 196.000 2528.700 ;
        RECT 4.000 2432.380 196.000 2527.540 ;
        RECT 4.000 2431.220 195.700 2432.380 ;
        RECT 4.000 2341.660 196.000 2431.220 ;
        RECT 4.300 2340.500 196.000 2341.660 ;
        RECT 4.000 2308.060 196.000 2340.500 ;
        RECT 4.000 2306.900 195.700 2308.060 ;
        RECT 4.000 2183.740 196.000 2306.900 ;
        RECT 4.000 2182.580 195.700 2183.740 ;
        RECT 4.000 2154.620 196.000 2182.580 ;
        RECT 4.300 2153.460 196.000 2154.620 ;
        RECT 4.000 2059.420 196.000 2153.460 ;
        RECT 4.000 2058.260 195.700 2059.420 ;
        RECT 4.000 1967.580 196.000 2058.260 ;
        RECT 4.300 1966.420 196.000 1967.580 ;
        RECT 4.000 1935.100 196.000 1966.420 ;
        RECT 4.000 1933.940 195.700 1935.100 ;
        RECT 4.000 1810.780 196.000 1933.940 ;
        RECT 4.000 1809.620 195.700 1810.780 ;
        RECT 4.000 1780.540 196.000 1809.620 ;
        RECT 4.300 1779.380 196.000 1780.540 ;
        RECT 4.000 1686.460 196.000 1779.380 ;
        RECT 4.000 1685.300 195.700 1686.460 ;
        RECT 4.000 1593.500 196.000 1685.300 ;
        RECT 4.300 1592.340 196.000 1593.500 ;
        RECT 4.000 1562.140 196.000 1592.340 ;
        RECT 4.000 1560.980 195.700 1562.140 ;
        RECT 4.000 1437.820 196.000 1560.980 ;
        RECT 4.000 1436.660 195.700 1437.820 ;
        RECT 4.000 1406.460 196.000 1436.660 ;
        RECT 4.300 1405.300 196.000 1406.460 ;
        RECT 4.000 1313.500 196.000 1405.300 ;
        RECT 4.000 1312.340 195.700 1313.500 ;
        RECT 4.000 1219.420 196.000 1312.340 ;
        RECT 4.300 1218.260 196.000 1219.420 ;
        RECT 4.000 1189.180 196.000 1218.260 ;
        RECT 4.000 1188.020 195.700 1189.180 ;
        RECT 4.000 1064.860 196.000 1188.020 ;
        RECT 4.000 1063.700 195.700 1064.860 ;
        RECT 4.000 1032.380 196.000 1063.700 ;
        RECT 4.300 1031.220 196.000 1032.380 ;
        RECT 4.000 940.540 196.000 1031.220 ;
        RECT 4.000 939.380 195.700 940.540 ;
        RECT 4.000 845.340 196.000 939.380 ;
        RECT 4.300 844.180 196.000 845.340 ;
        RECT 4.000 816.220 196.000 844.180 ;
        RECT 4.000 815.060 195.700 816.220 ;
        RECT 4.000 691.900 196.000 815.060 ;
        RECT 4.000 690.740 195.700 691.900 ;
        RECT 4.000 658.300 196.000 690.740 ;
        RECT 4.300 657.140 196.000 658.300 ;
        RECT 4.000 567.580 196.000 657.140 ;
        RECT 4.000 566.420 195.700 567.580 ;
        RECT 4.000 471.260 196.000 566.420 ;
        RECT 4.300 470.100 196.000 471.260 ;
        RECT 4.000 443.260 196.000 470.100 ;
        RECT 4.000 442.100 195.700 443.260 ;
        RECT 4.000 318.940 196.000 442.100 ;
        RECT 4.000 317.780 195.700 318.940 ;
        RECT 4.000 284.220 196.000 317.780 ;
        RECT 4.300 283.060 196.000 284.220 ;
        RECT 4.000 194.620 196.000 283.060 ;
        RECT 4.000 193.460 195.700 194.620 ;
        RECT 4.000 97.180 196.000 193.460 ;
        RECT 4.300 96.020 196.000 97.180 ;
        RECT 4.000 70.300 196.000 96.020 ;
        RECT 4.000 69.140 195.700 70.300 ;
        RECT 4.000 15.540 196.000 69.140 ;
      LAYER Metal4 ;
        RECT 82.460 20.810 98.740 1581.350 ;
        RECT 100.940 20.810 175.540 1581.350 ;
        RECT 177.740 20.810 191.380 1581.350 ;
  END
END user_proj_example
END LIBRARY

