VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 42.560 2800.000 43.120 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1280.160 4.000 1280.720 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1061.760 4.000 1062.320 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 843.360 4.000 843.920 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 624.960 4.000 625.520 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 406.560 4.000 407.120 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END io_in[15]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 260.960 2800.000 261.520 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 479.360 2800.000 479.920 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 697.760 2800.000 698.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 916.160 2800.000 916.720 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1134.560 2800.000 1135.120 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1352.960 2800.000 1353.520 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1571.360 2800.000 1571.920 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1716.960 4.000 1717.520 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1498.560 4.000 1499.120 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 188.160 2800.000 188.720 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1134.560 4.000 1135.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 916.160 4.000 916.720 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 697.760 4.000 698.320 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 479.360 4.000 479.920 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 4.000 261.520 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 4.000 43.120 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 406.560 2800.000 407.120 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 624.960 2800.000 625.520 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 843.360 2800.000 843.920 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1061.760 2800.000 1062.320 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1280.160 2800.000 1280.720 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1498.560 2800.000 1499.120 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1716.960 2800.000 1717.520 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1571.360 4.000 1571.920 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1352.960 4.000 1353.520 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 115.360 2800.000 115.920 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1207.360 4.000 1207.920 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 988.960 4.000 989.520 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 770.560 4.000 771.120 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 552.160 4.000 552.720 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 333.760 4.000 334.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END io_out[15]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 333.760 2800.000 334.320 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 552.160 2800.000 552.720 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 770.560 2800.000 771.120 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 988.960 2800.000 989.520 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1207.360 2800.000 1207.920 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1425.760 2800.000 1426.320 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1644.160 2800.000 1644.720 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1644.160 4.000 1644.720 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1425.760 4.000 1426.320 ;
    END
  END io_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 1740.780 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 1740.780 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 0.000 599.760 4.000 ;
    END
  END wb_rst_i
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1398.880 0.000 1399.440 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1798.720 0.000 1799.280 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2198.560 0.000 2199.120 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2598.400 0.000 2598.960 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 999.040 0.000 999.600 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 2793.280 1740.780 ;
      LAYER Metal2 ;
        RECT 8.540 4.300 2791.460 1740.670 ;
        RECT 8.540 4.000 199.060 4.300 ;
        RECT 200.220 4.000 598.900 4.300 ;
        RECT 600.060 4.000 998.740 4.300 ;
        RECT 999.900 4.000 1398.580 4.300 ;
        RECT 1399.740 4.000 1798.420 4.300 ;
        RECT 1799.580 4.000 2198.260 4.300 ;
        RECT 2199.420 4.000 2598.100 4.300 ;
        RECT 2599.260 4.000 2791.460 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1717.820 2796.000 1740.620 ;
        RECT 4.300 1716.660 2795.700 1717.820 ;
        RECT 4.000 1645.020 2796.000 1716.660 ;
        RECT 4.300 1643.860 2795.700 1645.020 ;
        RECT 4.000 1572.220 2796.000 1643.860 ;
        RECT 4.300 1571.060 2795.700 1572.220 ;
        RECT 4.000 1499.420 2796.000 1571.060 ;
        RECT 4.300 1498.260 2795.700 1499.420 ;
        RECT 4.000 1426.620 2796.000 1498.260 ;
        RECT 4.300 1425.460 2795.700 1426.620 ;
        RECT 4.000 1353.820 2796.000 1425.460 ;
        RECT 4.300 1352.660 2795.700 1353.820 ;
        RECT 4.000 1281.020 2796.000 1352.660 ;
        RECT 4.300 1279.860 2795.700 1281.020 ;
        RECT 4.000 1208.220 2796.000 1279.860 ;
        RECT 4.300 1207.060 2795.700 1208.220 ;
        RECT 4.000 1135.420 2796.000 1207.060 ;
        RECT 4.300 1134.260 2795.700 1135.420 ;
        RECT 4.000 1062.620 2796.000 1134.260 ;
        RECT 4.300 1061.460 2795.700 1062.620 ;
        RECT 4.000 989.820 2796.000 1061.460 ;
        RECT 4.300 988.660 2795.700 989.820 ;
        RECT 4.000 917.020 2796.000 988.660 ;
        RECT 4.300 915.860 2795.700 917.020 ;
        RECT 4.000 844.220 2796.000 915.860 ;
        RECT 4.300 843.060 2795.700 844.220 ;
        RECT 4.000 771.420 2796.000 843.060 ;
        RECT 4.300 770.260 2795.700 771.420 ;
        RECT 4.000 698.620 2796.000 770.260 ;
        RECT 4.300 697.460 2795.700 698.620 ;
        RECT 4.000 625.820 2796.000 697.460 ;
        RECT 4.300 624.660 2795.700 625.820 ;
        RECT 4.000 553.020 2796.000 624.660 ;
        RECT 4.300 551.860 2795.700 553.020 ;
        RECT 4.000 480.220 2796.000 551.860 ;
        RECT 4.300 479.060 2795.700 480.220 ;
        RECT 4.000 407.420 2796.000 479.060 ;
        RECT 4.300 406.260 2795.700 407.420 ;
        RECT 4.000 334.620 2796.000 406.260 ;
        RECT 4.300 333.460 2795.700 334.620 ;
        RECT 4.000 261.820 2796.000 333.460 ;
        RECT 4.300 260.660 2795.700 261.820 ;
        RECT 4.000 189.020 2796.000 260.660 ;
        RECT 4.300 187.860 2795.700 189.020 ;
        RECT 4.000 116.220 2796.000 187.860 ;
        RECT 4.300 115.060 2795.700 116.220 ;
        RECT 4.000 43.420 2796.000 115.060 ;
        RECT 4.300 42.260 2795.700 43.420 ;
        RECT 4.000 15.540 2796.000 42.260 ;
      LAYER Metal4 ;
        RECT 1096.060 533.210 1097.140 878.550 ;
        RECT 1099.340 533.210 1173.940 878.550 ;
        RECT 1176.140 533.210 1250.740 878.550 ;
        RECT 1252.940 533.210 1327.540 878.550 ;
        RECT 1329.740 533.210 1404.340 878.550 ;
        RECT 1406.540 533.210 1481.140 878.550 ;
        RECT 1483.340 533.210 1557.940 878.550 ;
        RECT 1560.140 533.210 1561.700 878.550 ;
  END
END user_proj_example
END LIBRARY

