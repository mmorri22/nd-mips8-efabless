magic
tech gf180mcuD
magscale 1 5
timestamp 1701656237
<< obsm1 >>
rect 672 1538 19320 298342
<< metal2 >>
rect 4928 0 4984 400
rect 14896 0 14952 400
<< obsm2 >>
rect 854 430 19418 298331
rect 854 400 4898 430
rect 5014 400 14866 430
rect 14982 400 19418 430
<< metal3 >>
rect 19600 292880 20000 292936
rect 0 290192 400 290248
rect 19600 280448 20000 280504
rect 0 271488 400 271544
rect 19600 268016 20000 268072
rect 19600 255584 20000 255640
rect 0 252784 400 252840
rect 19600 243152 20000 243208
rect 0 234080 400 234136
rect 19600 230720 20000 230776
rect 19600 218288 20000 218344
rect 0 215376 400 215432
rect 19600 205856 20000 205912
rect 0 196672 400 196728
rect 19600 193424 20000 193480
rect 19600 180992 20000 181048
rect 0 177968 400 178024
rect 19600 168560 20000 168616
rect 0 159264 400 159320
rect 19600 156128 20000 156184
rect 19600 143696 20000 143752
rect 0 140560 400 140616
rect 19600 131264 20000 131320
rect 0 121856 400 121912
rect 19600 118832 20000 118888
rect 19600 106400 20000 106456
rect 0 103152 400 103208
rect 19600 93968 20000 94024
rect 0 84448 400 84504
rect 19600 81536 20000 81592
rect 19600 69104 20000 69160
rect 0 65744 400 65800
rect 19600 56672 20000 56728
rect 0 47040 400 47096
rect 19600 44240 20000 44296
rect 19600 31808 20000 31864
rect 0 28336 400 28392
rect 19600 19376 20000 19432
rect 0 9632 400 9688
rect 19600 6944 20000 7000
<< obsm3 >>
rect 400 292966 19600 298326
rect 400 292850 19570 292966
rect 400 290278 19600 292850
rect 430 290162 19600 290278
rect 400 280534 19600 290162
rect 400 280418 19570 280534
rect 400 271574 19600 280418
rect 430 271458 19600 271574
rect 400 268102 19600 271458
rect 400 267986 19570 268102
rect 400 255670 19600 267986
rect 400 255554 19570 255670
rect 400 252870 19600 255554
rect 430 252754 19600 252870
rect 400 243238 19600 252754
rect 400 243122 19570 243238
rect 400 234166 19600 243122
rect 430 234050 19600 234166
rect 400 230806 19600 234050
rect 400 230690 19570 230806
rect 400 218374 19600 230690
rect 400 218258 19570 218374
rect 400 215462 19600 218258
rect 430 215346 19600 215462
rect 400 205942 19600 215346
rect 400 205826 19570 205942
rect 400 196758 19600 205826
rect 430 196642 19600 196758
rect 400 193510 19600 196642
rect 400 193394 19570 193510
rect 400 181078 19600 193394
rect 400 180962 19570 181078
rect 400 178054 19600 180962
rect 430 177938 19600 178054
rect 400 168646 19600 177938
rect 400 168530 19570 168646
rect 400 159350 19600 168530
rect 430 159234 19600 159350
rect 400 156214 19600 159234
rect 400 156098 19570 156214
rect 400 143782 19600 156098
rect 400 143666 19570 143782
rect 400 140646 19600 143666
rect 430 140530 19600 140646
rect 400 131350 19600 140530
rect 400 131234 19570 131350
rect 400 121942 19600 131234
rect 430 121826 19600 121942
rect 400 118918 19600 121826
rect 400 118802 19570 118918
rect 400 106486 19600 118802
rect 400 106370 19570 106486
rect 400 103238 19600 106370
rect 430 103122 19600 103238
rect 400 94054 19600 103122
rect 400 93938 19570 94054
rect 400 84534 19600 93938
rect 430 84418 19600 84534
rect 400 81622 19600 84418
rect 400 81506 19570 81622
rect 400 69190 19600 81506
rect 400 69074 19570 69190
rect 400 65830 19600 69074
rect 430 65714 19600 65830
rect 400 56758 19600 65714
rect 400 56642 19570 56758
rect 400 47126 19600 56642
rect 430 47010 19600 47126
rect 400 44326 19600 47010
rect 400 44210 19570 44326
rect 400 31894 19600 44210
rect 400 31778 19570 31894
rect 400 28422 19600 31778
rect 430 28306 19600 28422
rect 400 19462 19600 28306
rect 400 19346 19570 19462
rect 400 9718 19600 19346
rect 430 9602 19600 9718
rect 400 7030 19600 9602
rect 400 6914 19570 7030
rect 400 1554 19600 6914
<< metal4 >>
rect 2224 1538 2384 298342
rect 9904 1538 10064 298342
rect 17584 1538 17744 298342
<< obsm4 >>
rect 8246 2081 9874 158135
rect 10094 2081 17554 158135
rect 17774 2081 19138 158135
<< labels >>
rlabel metal3 s 19600 6944 20000 7000 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 19600 44240 20000 44296 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 19600 81536 20000 81592 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 19600 118832 20000 118888 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 19600 156128 20000 156184 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 19600 193424 20000 193480 6 io_in[5]
port 6 nsew signal input
rlabel metal3 s 19600 230720 20000 230776 6 io_in[6]
port 7 nsew signal input
rlabel metal3 s 19600 268016 20000 268072 6 io_in[7]
port 8 nsew signal input
rlabel metal3 s 19600 31808 20000 31864 6 io_oeb[0]
port 9 nsew signal output
rlabel metal3 s 0 196672 400 196728 6 io_oeb[10]
port 10 nsew signal output
rlabel metal3 s 0 159264 400 159320 6 io_oeb[11]
port 11 nsew signal output
rlabel metal3 s 0 121856 400 121912 6 io_oeb[12]
port 12 nsew signal output
rlabel metal3 s 0 84448 400 84504 6 io_oeb[13]
port 13 nsew signal output
rlabel metal3 s 0 47040 400 47096 6 io_oeb[14]
port 14 nsew signal output
rlabel metal3 s 0 9632 400 9688 6 io_oeb[15]
port 15 nsew signal output
rlabel metal3 s 19600 69104 20000 69160 6 io_oeb[1]
port 16 nsew signal output
rlabel metal3 s 19600 106400 20000 106456 6 io_oeb[2]
port 17 nsew signal output
rlabel metal3 s 19600 143696 20000 143752 6 io_oeb[3]
port 18 nsew signal output
rlabel metal3 s 19600 180992 20000 181048 6 io_oeb[4]
port 19 nsew signal output
rlabel metal3 s 19600 218288 20000 218344 6 io_oeb[5]
port 20 nsew signal output
rlabel metal3 s 19600 255584 20000 255640 6 io_oeb[6]
port 21 nsew signal output
rlabel metal3 s 19600 292880 20000 292936 6 io_oeb[7]
port 22 nsew signal output
rlabel metal3 s 0 271488 400 271544 6 io_oeb[8]
port 23 nsew signal output
rlabel metal3 s 0 234080 400 234136 6 io_oeb[9]
port 24 nsew signal output
rlabel metal3 s 19600 19376 20000 19432 6 io_out[0]
port 25 nsew signal output
rlabel metal3 s 0 215376 400 215432 6 io_out[10]
port 26 nsew signal output
rlabel metal3 s 0 177968 400 178024 6 io_out[11]
port 27 nsew signal output
rlabel metal3 s 0 140560 400 140616 6 io_out[12]
port 28 nsew signal output
rlabel metal3 s 0 103152 400 103208 6 io_out[13]
port 29 nsew signal output
rlabel metal3 s 0 65744 400 65800 6 io_out[14]
port 30 nsew signal output
rlabel metal3 s 0 28336 400 28392 6 io_out[15]
port 31 nsew signal output
rlabel metal3 s 19600 56672 20000 56728 6 io_out[1]
port 32 nsew signal output
rlabel metal3 s 19600 93968 20000 94024 6 io_out[2]
port 33 nsew signal output
rlabel metal3 s 19600 131264 20000 131320 6 io_out[3]
port 34 nsew signal output
rlabel metal3 s 19600 168560 20000 168616 6 io_out[4]
port 35 nsew signal output
rlabel metal3 s 19600 205856 20000 205912 6 io_out[5]
port 36 nsew signal output
rlabel metal3 s 19600 243152 20000 243208 6 io_out[6]
port 37 nsew signal output
rlabel metal3 s 19600 280448 20000 280504 6 io_out[7]
port 38 nsew signal output
rlabel metal3 s 0 290192 400 290248 6 io_out[8]
port 39 nsew signal output
rlabel metal3 s 0 252784 400 252840 6 io_out[9]
port 40 nsew signal output
rlabel metal4 s 2224 1538 2384 298342 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 298342 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 298342 6 vss
port 42 nsew ground bidirectional
rlabel metal2 s 4928 0 4984 400 6 wb_clk_i
port 43 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 wb_rst_i
port 44 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3976274
string GDS_FILE /mnt/c/Users/mmorri22/caravel_user_project/openlane/user_proj_example/runs/23_12_03_21_15/results/signoff/user_proj_example.magic.gds
string GDS_START 335636
<< end >>

